module dff (
    clock,
    reset,
    d_in,
    Q_out,
    Qb_out
);

  //Step1 : Declare Port Directions
  input clock, reset, d_in;
  output reg Q_out, Qb_out;

  /*Understand the Behaviour of D flip-flop &
   check the coding style of synchronous reset*/

  always @(posedge clock) begin
    if (reset) Q_out <= 1'b0;
    else Q_out <= d_in;
  end

  //Step2 : Write the logic for Qbar	
  always @(posedge clock) begin
    if (reset) Qb_out <= 1'b1;
    else Qb_out <= ~d_in;
  end

endmodule
